module gi

pub struct Typelib {
	c &C.GITypelib
}
