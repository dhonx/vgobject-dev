module main

import gi

fn main() {
	repo := gi.Repository{}
	// repo.require('Gtk', '', .lazy)
	
	// n_infos := repo.get_n_infos('Gtk')
	// println(n_infos)

	// a := C.GI_FIELD_IS_READABLE

	// loaded_ns := repo.get_loaded_namespaces()
	// println(loaded_ns)
}
